module KeyBoard (input wire a, output reg b);



endmodule